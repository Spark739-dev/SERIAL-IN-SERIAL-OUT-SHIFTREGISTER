library verilog;
use verilog.vl_types.all;
entity siso_vlg_vec_tst is
end siso_vlg_vec_tst;
